* Rheostat, 2ohm total resistance

.subckt Rheostat left right up rsum=999k
B1 left  up I=V(left ,up)/(rsum*V(v_r))
B2 right up I=V(right,up)/(rsum*(1-V(v_r)))
.ends
